BRAKEREG.CIR - LINEAR ACTUATOR EXTERNAL CURRENT REGULATOR
.MODEL 2n6288 npn
+IS=7.86858e-13 BF=455.929 NF=0.85 VAF=10
+IKF=0.902779 ISE=2.00343e-13 NE=1.96023 BR=28.7722
+NR=1.5 VAR=1.12144 IKR=9.02779 ISC=4.92338e-16
+NC=3.9992 RB=8.77246 IRB=0.1 RBM=0.1
+RE=0.0001 RC=0.416835 XTB=0.1 XTI=2.87011
+EG=1.206 CJE=1.84157e-10 VJE=0.99 MJE=0.347174
+TF=7.13242e-09 XTF=1.50205 VTF=1.00686 ITF=0.998053
+CJC=1.06717e-10 VJC=0.942695 MJC=0.245406 XCJC=0.8
+FC=0.53342 CJS=0 VJS=0.75 MJS=0.5
+TR=2.97071e-08 PTF=0 KF=0 AF=1
* Model generated on Jan 24, 2004
* Model format: SPICE3
*
V_1	1	2	SIN(0 1 10)
V_2	9	0	DC	12
*
R_1	1	3	2
R_2	8	9	1
*
Q_1	2	2	4	2n6288
Q_2	3	3	4	2n6288
Q_3	7	7	2	2n6288
Q_4	7	7	3	2n6288
Q_5	4	4	5	2n6288
Q_6	5	6	7	2n6288
Q_7	8	4	6	2n6288
Q_8	6	6	0	2n6288
*
.IC	V(1)=0 V(2)=0 V(3)=0 V(4)=0 V(5)=0 V(6)=0 V(7)=0 V(8)=0
.TRAN	.001	.2	UIC
*
.PLOT	TRAN	V_1#branch V_2#branch
